library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity arccos_calculator is
	port (
		clk 	: in std_logic;
		reset : in std_logic;
		X 		: in std_logic_vector(7 downto 0);
		ANGLE : out std_logic_vector(9 downto 0)
	);
end arccos_calculator;

architecture rtl of arccos_calculator is
	signal X_i 	: SIGNED (7 downto 0);
	signal X2 	: SIGNED (15 downto 0);
	signal P1 	: SIGNED (6 downto 0);
	signal P2 	: SIGNED (8 downto 0);
	signal P3 	: SIGNED (8 downto 0);
	signal S1 	: SIGNED (8 downto 0);
	signal S2 	: SIGNED (10 downto 0);

begin
	-- X2 = X*X
	X2 <= X_i*X_i;
			
	-- P1 = (86*X2)/2^16
	P1 <= resize(shift_right((to_signed(86, 8)*X2), 16), 7);
	
	-- S1 = 191 + P1
	S1 <= resize(to_signed(191, 8) + P1, 9);
	
	-- P2 = (S1*X2)/2^16
	P2 <= resize(shift_right((S1*X2), 16), 9);

	-- S2 = 1144 + P2
	S2 <= to_signed(1144, 11) + P2;
	
	-- P3 = (S2*X)/2^9
	P3 <= resize(shift_right((S2*signed(X_i)), 9), 9);
	
	calculate_angle : process (clk, reset)
		
	begin
		if (reset = '1') then
			ANGLE <= (others => '0');
			X_i <= (others => '0');
		elsif (rising_edge(clk)) then
			X_i <= signed(X);
			
			-- ANGLE = 900 - P3
			ANGLE <= std_logic_vector((to_signed(900, 10) - P3));
		end if;
	end process calculate_angle;
end rtl;